# ====================================================================
#
#      gpio.cdl
#
#      Generic API for accessing GPIO
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008, 2009 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
#    
# Contributors:
# Date:           2010-10-23
#
#####DESCRIPTIONEND####
# ====================================================================

cdl_package CYGPKG_IO_GPIO {

    display    "Generic API definition for accessing GPIO"
    
    requires    CYGINT_IO_GPIO_ROUTINE

    include_dir "cyg/io/"
    
    description "
        The GPIO package provides generic definitions to access and
        configure the General Purpose IOs."

    cdl_interface CYGINT_IO_GPIO_ROUTINE {
    display   "HAL supports GPIO access."
    description "
          The IO GPIO package provides the GPIO access definition headers.
          The actual GPIO routines are to be implemented on HAL bases."
    }

}
