# ==========================================================================
#
#      stm32_r6_fb.cdl
#
#      r61523 LCD controller platform specific code
#
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2014 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    ccoutand
# Contributors: 
# Date:         2011-07-01
# Purpose:      
# Description:  r61523 LCD controller platform specific code (STM32 R6)
#
#####DESCRIPTIONEND####
#
# ===========================================================================

cdl_package CYGPKG_DEVS_FRAMEBUF_CORTEXM_STM32_R6 {
    display       "Platform specific device driver for r61523 LCD controller ((STM32 R6)"
    parent        CYGPKG_DEVS_FRAMEBUF_R61523
    active_if     CYGPKG_IO_FRAMEBUF
    active_if     CYGPKG_DEVS_FRAMEBUF_R61523
    active_if     CYGPKG_HAL_CORTEXM_STM32

    implements    CYGINT_DEVS_FRAMEBUF_R61523_PLF

    include_dir   cyg/io
    compile       r61523_plf.c

    description   "
        This package provides the macros necessary for the r61523 
        framebuffer device driver to access the hardware. The r61523
        LCD controller initialization sequence is also provided by 
        this package."

    define_proc {
        puts $::cdl_system_header "#define CYGPKG_DEVS_FRAMEBUF_R61523_PLF_H <pkgconf/devs_framebuf_cortexm_stm32_r6.h>"
        puts $::cdl_system_header "#define CYGPKG_DEVS_FRAMEBUF_R61523_PLF_INL <cyg/io/r61523_plf.inl>"
    }

    cdl_component CYGPKG_DEVS_FRAMEBUF_CORTEXM_STM32_R6_OPTIONS {
        display       "STM32 R6 Framebuffer build options"
        flavor        none
        description   "
            Package specific build options including control over
            compiler flags used only in building the generic frame
            buffer package, and details of which tests are built."

        cdl_option CYGPKG_DEVS_FRAMEBUF_CORTEXM_STM32_R6_TESTS {
            display      "STM32 R6 Framebuffer tests"
            active_if    CYGINT_IO_FRAMEBUF_DEVICES
            flavor       data
            calculated   { "tests/stm32_r6_fb" }
            description "
                This option specifies the set of tests for the STM32 R6 framebuffer package"
        }
    }
}