# ====================================================================
#
#      flash_mini_stm32.cdl
#
#      FLASH memory - Hardware support on MINI STM32 board
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
# Original data:  gthomas
# Contributors:   gthomas
# Date:           2011-05-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_CORTEXM_MINI_STM32 {
    display       "MINI STM32 FLASH memory support"
    description   "Hardware support on MINI STM32 board"

    parent        CYGPKG_IO_FLASH
    active_if     CYGPKG_IO_FLASH
    requires      CYGPKG_HAL_CORTEXM_STM32
    requires      CYGHWR_DEVS_SPI_CORTEXM_STM32_BUS1

    compile       -library=libextras.a flash_mini_stm32.c

    cdl_option CYGPKG_DEVS_FLASH_CORTEXM_MINI_STM32_TESTS {
        display     "Mini STM32 SPI Flash tests"
        active_if    CYGPKG_KERNEL
        active_if    CYGPKG_IO_SPI
        flavor       data
        no_define
        calculated { "tests/flash_mini_stm32_test" }
        description   "
            This option specifies the set of tests for the
            Mini STM32 SPI Flash."
    }
}

# EOF flash_mini_stm32.cdl
