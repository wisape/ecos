# ====================================================================
#
#      pwm_stm32.cdl
#
#      eCos STM32 PWM configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2010 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Wisape <wisape@gmail.com>
# Contributors:
# Date:           2015-06-14
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_PWM_CORTEXM_STM32 {
    display     "PWM bus driver for STM32 family of CortexM controllers"
    
    parent      CYGPKG_IO
    active_if   CYGPKG_IO
    active_if   CYGPKG_HAL_CORTEXM_STM32 

    description " 
           This package provides a generic PWM device driver for the on-chip
           PWM peripherals in STM32 processors."
           
    include_dir cyg/io
    compile     pwm_stm32.c

    define_proc {
      puts $::cdl_system_header "#define CYGDAT_DEVS_STM32_PWM_INL <cyg/io/pwm_stm32.inl>"
    }

    cdl_option CYGDAT_DEVS_STM32_PWM_NAME {
        display "Device name for stm32 pwm"

        flavor data

        default_value {"\"/dev/pwm\""}

        description "The package specifies the name of stm32 pwm."
    }
    
}
