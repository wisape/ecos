# ====================================================================
#
#      libpng.cdl
#
#      libpng is the official PNG reference library
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2014 Free Software Foundation, Inc.                  
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
# Original data:  http://www.libpng.org/pub/png/libpng.html
#                 Version:
#                 1.6.10rc1
# Contributors:
# Date:           2014-05-29
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_LIBPNG {
    display     "PNG graphical library"
    requires    CYGPKG_LIBC_STDIO
    requires    CYGPKG_LIBC_STDLIB
    requires    CYGPKG_LIBC_STRING
    requires    CYGPKG_LIBC_SETJMP
    requires    CYGPKG_ISOINFRA
    requires    CYGPKG_MEMALLOC
    requires    CYGPKG_COMPRESS_ZLIB
    requires    CYGPKG_CRC

    include_dir cyg/libpng

    compile png.c pngerror.c pngget.c pngmem.c pngpread.c pngread.c pngrio.c 
    compile pngrtran.c pngrutil.c pngset.c pngtrans.c pngwio.c pngwrite.c 
    compile pngwtran.c pngwutil.c

    description "
        This package includes support for the libPNG 1.6.11rc1"

    cdl_component CYGPKG_LIBPNG_OPTIONS {
        display       "libPNG library build options"
        flavor        none
        description   "
        Package specific build options including control over
        compiler flags used only in building this package,
        and details of which tests are built."

        cdl_option CYGPKG_LIBPNG_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D__ECOS__" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_LIBPNG_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this package. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGTST_LIBPNG_BUILD_TESTS {
        display       "Build LibPNG tests"
        flavor         bool
        no_define
        default_value  0
        active_if      CYGPKG_FS_ROM_TESTS
        active_if      CYGINT_IO_FRAMEBUF_DEVICES

        cdl_option CYGPKG_LIBPNG_TESTS {
            display    "LibPNG tests"
            flavor      data
            no_define
            calculated { "tests/readpng" }
            description   "
                This option specifies the set of tests for the LibPNG 
                package."
        }
    }

}
