# ====================================================================
#
#      mb_uart_lite.cdl
#
#      Microblaze UART Lite serial configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
# Original data:  
# Contributors:
# Date:           2011-03-05
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_IO_SERIAL_MICROBLAZE_UARTLITE {
    display       "Microblaze UART Lite serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL
    active_if     CYGPKG_HAL_MICROBLAZE

    compile       -library=libextras.a  mb_uart_lite.c

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_DEVICE_HEADER <pkgconf/io_serial_microblaze_uartlite.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_SERIAL_A {
    display       "Microblaze serial port A driver"
    flavor        bool
    default_value 1
    requires      (CYGIMP_KERNEL_INTERRUPTS_CHAIN || \
                      !CYGPKG_IO_SERIAL_MICROBLAZE_SERIAL_B)
    description   "
        This option includes the serial device driver for the Microblaze 
        port A. If both drivers need to be enabled, interrupt
        chaining must be enabled in the kernel configuration."

    cdl_option CYGDAT_IO_SERIAL_MICROBLAZE_SERIAL_A_NAME {
        display       "Device name for the Microblaze serial port A"
        flavor        data
        default_value {"\"/dev/ser0\""}
        description   "
            This option specifies the device name for the Microblaze
            port A."
    }

    cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_SERIAL_A_BUFSIZE {
        display       "Buffer size for the Microblaze serial port A driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used for 
            the Microblaze port A."
    }

    cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_SERIAL_A_IOBASE {
        display       "I/O base address for the Microblaze serial port 0"
        flavor        data
        default_value 0x8F800000
            description "
            This option specifies the I/O address of for the serial port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_SERIAL_A_INT {
        display        "INT for the Microblaze serial port 0"
        flavor         data
        default_value  3
        legal_values   0 to CYGNUM_HAL_MICROBLAZE_IPC_MAXIRQ
            description "
            This option specifies the interrupt vector for the serial port 0."
    }
}
cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_SERIAL_B {
    display       "Microblaze serial port B driver"
    flavor        bool
    default_value 0
    description   "
        This option includes the serial device driver for the Microblaze
        port B."

    cdl_option CYGDAT_IO_SERIAL_MICROBLAZE_SERIAL_B_NAME {
        display       "Device name for the Microblaze serial port B"
        flavor        data
        default_value {"\"/dev/ser1\""}
        description   "
            This option specifies the device name for the Microblaze
            port B."
    }

    cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_SERIAL_B_BUFSIZE {
        display       "Buffer size for the Microblaze serial port B driver"
        flavor        data
        legal_values  0 to 8192
        default_value 128
        description   "
            This option specifies the size of the internal buffers used 
            for the Microblaze port B."
    }

    cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_SERIAL_B_IOBASE {
        display       "I/O base address for the Microblaze serial port 0"
        flavor        data
        default_value 0x8F800000
            description "
            This option specifies the I/O address of for the serial port 0."
    }

    cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_SERIAL_B_INT {
        display        "INT for the Microblaze serial port 0"
        flavor         data
        default_value  3
        legal_values   0 to CYGNUM_HAL_MICROBLAZE_IPC_MAXIRQ
            description "
            This option specifies the interrupt vector for the serial port 0."
    }
}

    cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
        Package specific build options including control over
        compiler flags used only in building this package,
        and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_MICROBLAZE_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_MICROBLAZE_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_MICROBLAZE_SERIAL_B

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_MICROBLAZE_SERIAL_B_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"microblaze\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF mb_uart_lite.cdl
