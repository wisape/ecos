# ====================================================================
#
#      mb_uart16550.cdl
#
#      eCos serial PC configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      ccoutand
# Original data:  i386
# Contributors:   jskov
# Date:           2011-02-18
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_IO_SERIAL_MICROBLAZE_UART16550 {
    display       "Microblaze serial device drivers"

    parent        CYGPKG_IO_SERIAL_DEVICES
    active_if     CYGPKG_IO_SERIAL

    requires      CYGPKG_ERROR
    requires      CYGPKG_IO_SERIAL_GENERIC_16X5X
    include_dir   cyg/io
    description   "
           This option enables the serial device drivers for the PC."

    # FIXME: This really belongs in the GENERIC_16X5X package
    cdl_interface CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED {
        display   "Generic 16x5x serial driver required"
    }
    define_proc {
        puts $::cdl_header "#define CYGPRI_IO_SERIAL_GENERIC_16X5X_STEP 4"
    }

    define_proc {
        puts $::cdl_system_header "/***** serial driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_INL <cyg/io/mb_uart16550.inl>"
        puts $::cdl_system_header "#define CYGDAT_IO_SERIAL_GENERIC_16X5X_CFG <pkgconf/io_serial_microblaze_uart16550.h>"
        puts $::cdl_system_header "/*****  serial driver proc output end  *****/"
    }

    cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0 {
        display       "Microblaze serial port 0 driver"
        flavor        bool
        default_value 1
        description   "
            This option includes the serial device driver for port 0 on the 
            Microblaze."

        implements    CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
        implements    CYGINT_IO_SERIAL_FLOW_CONTROL_HW
        implements    CYGINT_IO_SERIAL_LINE_STATUS_HW

        cdl_option CYGDAT_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0_NAME {
            display       "Device name for Microblaze serial port 0"
            flavor        data
            default_value {"\"/dev/ser0\""}
            description   "
                This option specifies the device name port 0 on the Microblaze."
        }

        cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0_BAUD {
            display       "Baud rate for the Microblaze serial port 0 driver"
            flavor        data
            legal_values  { 3600 4800 9600 38400 57600 115200 }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed) for the
                Microblaze port 0."
        }

        cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0_BUFSIZE {
            display       "Buffer size for the Microblaze serial port 0 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used
                for the Microblaze port 0."
        }

        cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0_IOBASE {
            display "I/O base address for the Microblaze serial port 0"
            flavor    data
            default_value 0x8F800000
            description "
            This option specifies the I/O address of the 16550 for serial port 0."
        }

       cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0_INT {
            display        "INT for the Microblaze serial port 0"
            flavor         data
            default_value  3
            legal_values   0 to CYGNUM_HAL_MICROBLAZE_IPC_MAXIRQ
            description "
            This option specifies the interrupt vector of the 16550 for serial port 0."
       }

       cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0_CLKFREQ {
            display        "Clock frequency for the Microblaze serial port 0"
            flavor          data
            default_value   { CYGNUM_HAL_MICROBLAZE_SYSCLOCK_FREQ }
            description "
            This option specifies the clock frequency of the 16550 for serial port 0."
       }
    }

    cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_UART16550_SERIAL1 {
        display       "Microblaze serial port 1 driver"
        flavor        bool
        default_value 0
        description   "
            This option includes the serial device driver for port 1 on
            the Microblaze."

        implements    CYGINT_IO_SERIAL_GENERIC_16X5X_REQUIRED
        implements    CYGINT_IO_SERIAL_FLOW_CONTROL_HW
        implements    CYGINT_IO_SERIAL_LINE_STATUS_HW

        cdl_option CYGDAT_IO_SERIAL_MICROBLAZE_UART16550_SERIAL1_NAME {
            display       "Device name for Microblaze serial port 1"
            flavor        data
            default_value {"\"/dev/ser1\""}
            description   "
                This option specifies the device name port 1 on the Microblaze."
        }

        cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL1_BAUD {
            display       "Baud rate for the Microblaze serial port 1 driver"
            flavor        data
            legal_values  { 3600 4800 9600 38400 57600 115200 }
            default_value 38400
            description   "
                This option specifies the default baud rate (speed) for the
                Microblaze port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL1_BUFSIZE {
            display       "Buffer size for the Microblaze serial port 1 driver"
            flavor        data
            legal_values  0 to 8192
            default_value 128
            description   "
                This option specifies the size of the internal buffers used
                for the Microblaze port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL1_IOBASE {
            display "I/O base address for the Microblaze serial port 1"
            flavor    data
            default_value 0x8F800000
            description "
            This option specifies the I/O address of the 16550 for serial port 1."
        }

        cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL1_INT {
            display       "INT for the Microblaze serial port 1"
            flavor         data
            default_value  3
            legal_values   0 to CYGNUM_HAL_MICROBLAZE_IPC_MAXIRQ
            description "
            This option specifies the interrupt vector of the 16550 for serial port 1."
        }

       cdl_option CYGNUM_IO_SERIAL_MICROBLAZE_UART16550_SERIAL1_CLKFREQ {
            display        "Clock frequency for the Microblaze serial port "
            flavor          data
            default_value   { CYGNUM_HAL_MICROBLAZE_SYSCLOCK_FREQ }
            description "
            This option specifies the clock frequency of the 16550 for serial port 1."
       }
    }

    cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_UART16550_OPTIONS {
        display "Serial device driver build options"
        flavor  none
        description   "
        Package specific build options including control over
        compiler flags used only in building this package,
        and details of which tests are built."


        cdl_option CYGPKG_IO_SERIAL_MICROBLAZE_UART16550_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_IO_SERIAL_MICROBLAZE_UART16550_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGPKG_IO_SERIAL_MICROBLAZE_UART16550_TESTING {
        display    "Testing parameters"
        flavor     bool
        calculated 1
        active_if  CYGPKG_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0

        cdl_option CYGPRI_SER_TEST_SER_DEV {
            display       "Serial device used for testing"
            flavor        data
            default_value { CYGDAT_IO_SERIAL_MICROBLAZE_UART16550_SERIAL0_NAME }
        }

        define_proc {
            puts $::cdl_header "#define CYGPRI_SER_TEST_CRASH_ID \"Microblaze\""
            puts $::cdl_header "#define CYGPRI_SER_TEST_TTY_DEV  \"/dev/tty0\""
        }
    }
}

# EOF mb_uart16550.cdl
