#==========================================================================
#
#      hal_freescale_qman.cdl
#
#      Freescale DPAA Queue Manager
#
#==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                           
## -------------------------------------------                             
## This file is part of eCos, the Embedded Configurable Operating System.  
## Copyright (C) 2013 Free Software Foundation, Inc.                       
##
## eCos is free software; you can redistribute it and/or modify it under   
## the terms of the GNU General Public License as published by the Free    
## Software Foundation; either version 2 or (at your option) any later     
## version.                                                                
##
## eCos is distributed in the hope that it will be useful, but WITHOUT     
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or   
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License   
## for more details.                                                       
##
## You should have received a copy of the GNU General Public License       
## along with eCos; if not, write to the Free Software Foundation, Inc.,   
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.           
##
## As a special exception, if other files instantiate templates or use     
## macros or inline functions from this file, or you compile this file     
## and link it with other works to produce a work based on this file,      
## this file does not by itself cause the resulting work to be covered by  
## the GNU General Public License. However the source code for this file   
## must still be made available in accordance with section (3) of the GNU  
## General Public License v2.                                              
##
## This exception does not invalidate any other reasons why a work based   
## on this file might be covered by the GNU General Public License.        
## -------------------------------------------                             
## ####ECOSGPLCOPYRIGHTEND####                                             
#==========================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    ccoutand
# Contributors:
# Date:         2013-01-21
#
#####DESCRIPTIONEND####
#
#==========================================================================
cdl_package CYGPKG_HAL_POWERPC_FREESCALE_DPAA_QMAN {
    display       "Freescale DPAA Queue Manager Interface"

    parent        CYGPKG_HAL_POWERPC
    active_if     CYGPKG_HAL_POWERPC_QORIQ_E500MC
    requires      CYGPKG_HAL_POWERPC_FREESCALE_DPAA_BMAN
    requires      CYGPKG_HAL_POWERPC_FREESCALE_DPAA_FMAN
    requires      CYGPKG_CRC
    include_dir   cyg/io

    description   "Queue Manager device driver for QoriQ processor"
    compile       -library=libextras.a fman.c

    cdl_option CYGPKG_HAL_POWERPC_FREESCALE_DPAA_QMAN_CHATTER {
        display         "Display status messages during FMAN operations"
        flavor           bool
        default_value    0
        description     "
           Selecting this option will cause the QMAN code to print status
           messages as various Ethernet operations are undertaken."
    }

    cdl_component CYGPKG_HAL_POWERPC_FREESCALE_DPAA_QMAN_OPTIONS {
        display  "Freescale Frame Manager driver build options"
        flavor   none
        no_define

        cdl_option CYGPKG_HAL_POWERPC_FREESCALE_DPAA_QMAN_CFLAGS_ADD {
            display       "Additional compiler flags"
            flavor         data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the frame manager driver package. 
                These flags are used in addition to the set of global 
                flags."
        }

        cdl_option CYGPKG_HAL_POWERPC_FREESCALE_DPAA_QMAN_CFLAGS_REMOVE {
            display        "Suppressed compiler flags"
            flavor         data
            no_define
            default_value { "" }
            description    "
                This option modifies the set of compiler flags for
                building the frame manager driver package. These flags 
                are removed from the set of global flags if present."
        }
    }

}