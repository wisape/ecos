# ====================================================================
#
#      nrf24l01.cdl
#
#      eCos 2.4G RF nrf24l01 configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      wisape
# Contributors:   
# Date:           2015-08-05
#
#####DESCRIPTIONEND####
#
# ====================================================================


cdl_package CYGPKG_DEVS_COMM_SPI_NRF24L01 {
    display     "NRF24L01 hardware interface"
    
    requires    CYGPKG_IO_SPI
    
    description " 
           This package provides 2.4G RF nrf24l01 interface."
           
    include_dir cyg/io
    
    compile  -library=libextras.a nrf24l01.c

    define_proc {
      puts $::cdl_system_header "#define CYGDAT_DEVS_NRF24L01_INL <cyg/io/nrf24l01.inl>"
    }
    
    cdl_option CYGDAT_DEVS_COMM_NRF24L01_NAME {
        display "Device name for 2.4G RF nrf24l01"

        flavor data

        default_value {"\"/dev/nrf24l01\""}

        description "The package specifies the name of 2.4G RF nrf24l01."
    }
}
