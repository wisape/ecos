# ==========================================================================
#
#      hal_powerpc_mpc8572ds.cdl
#
#      Freescale MPC8572DS evaluation board (MPC8572)
#
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    ccoutand
# Contributors: 
# Date:         2009-11-01
# Purpose:      
# Description:  HAL package configuration data
#
#####DESCRIPTIONEND####
#
# ==========================================================================

cdl_package CYGPKG_HAL_POWERPC_MPC8572DS {
    display       "Freescale MPC8572DS evaluation board "
    parent        CYGPKG_HAL_POWERPC
    requires      CYGPKG_HAL_POWERPC_QUICC3
    requires     ( CYGHWR_HAL_POWERPC_QUICC3=="MPC8572E" )

    define_header hal_powerpc_mpc8572ds.h
    include_dir   cyg/hal
    description   "
        The MPC8572DS HAL package provides the support needed to run
        eCos on a Freescale MPC8572DS evaluation board."

    compile       hal_diag.c hal_aux.c mpc8572ds.S plf_misc.c

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_PROFILE_HAL_TIMER
    requires      CYGSEM_HAL_POWERPC_RESET_USES_JUMP

    requires      { is_active(CYGPKG_DEVS_ETH_PHY) implies
                    (1 == CYGHWR_DEVS_ETH_PHY_VSC8244) }

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_powerpc_quicc3.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_powerpc_mpc8572ds.h>"

        puts $::cdl_header "#define HAL_PLATFORM_CPU  \"PowerPC MPC8572\""
        puts $::cdl_header "#define HAL_PLATFORM_BOARD \"MPC8572DS \""
        puts $::cdl_header "#define HAL_PLATFORM_EXTRA  \"\""
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  { "RAM" "ROM" "ROMRAM" }
        default_value { "RAM" }
    no_define
    define -file system.h CYG_HAL_STARTUP
        description   "
           This option is used to control where the application program will
           run, either from RAM or ROM (flash) memory.  ROM based applications
           must be self contained, while RAM applications will typically assume
           the existence of a debug environment, such as GDB stubs."
    }

    cdl_option CYGHWR_HAL_POWERPC_DISABLE_MMU {
        display       "DISABLE MMU"
        flavor        bool
        default_value 0
        description   "
            This option will disable the MMU enabled."
    }

    cdl_option CYGHWR_HAL_POWERPC_MPC8572DS_DDR1_CONTROLLER {
        display       "Configure DDR1 memory controller"
        flavor        bool
        default_value 1
        description   "
            Enable this option to configure the DDR1 memory controller"
    }

    cdl_option CYGHWR_HAL_POWERPC_MPC8572DS_DDR2_CONTROLLER {
        display       "Configure DDR2 memory controller"
        flavor        bool
        default_value 1
        requires { (CYGHWR_HAL_POWERPC_MPC8572DS_DDR1_CONTROLLER == 1) }
        description   "
            Enable this option to configure the DDR2 memory controller. Current 
            implementation does not allow to use DDR2 controller without DDR1 
            controller, some registers must be adjusted in that case (CS0_BNDS etc..)"
    }

     cdl_option CYGHWR_HAL_POWERPC_MPC8572DS_DDR_INTERLEAVED {
        display       "Configure DDR memory in interleaved mode"
        flavor        bool
        default_value 1
        description   "
            Enable this option to configure the DDR memory controller in interleaved mode."
    }

    cdl_option CYGHWR_HAL_POWERPC_MPC8572DS_SYS_CLK {
        display          "System Clock (MHz)"
        flavor           data
        default_value    100
        description      "
            MPC8572DS evaluation board system clock frequency in MHz (input clock)"
    }

    cdl_option CYGHWR_HAL_POWERPC_MPC8572DS_SYS_CLK_RATIO {
        display          "System Clock Ratio"
        flavor           data
        default_value    6
        legal_values     {4 5 6 8 10 12}
        description      "
            MPC8572DS evaluation board system clock ration (cfg_sys_pll)"
    }

    cdl_option CYGHWR_HAL_POWERPC_CPU_SPEED {
        display          "CPU CCB clock frequency (MHz)"
        flavor           data
        calculated       { CYGHWR_HAL_POWERPC_MPC8572DS_SYS_CLK * CYGHWR_HAL_POWERPC_MPC8572DS_SYS_CLK_RATIO }
        description      "
            MPC8572DS evaluation board CCB clock runs at 600MHz. This is the default setting, 
            with SYS_CLK configured to 100MHz and CFG_SYS_PLL set to 6."
    }

    cdl_option CYGHWR_HAL_POWERPC_MPC8572DS_CORE0_PLL_RATIO {
        display          "Core0 PLL Ration"
        flavor           data
        default_value    2.5
        legal_values     {1.5 2 2.5 3 3.5}
        description      "
            MPC8572DS evaluation board core0 PLL ratio (cfg_core0_pll)"
    }

    cdl_option CYGHWR_HAL_POWERPC_MPC8572DS_CORE1_PLL_RATIO {
        display          "Core1 PLL Ration"
        flavor           data
        default_value    2.5
        legal_values     {1.5 2 2.5 3 3.5}
        description      "
            MPC8572DS evaluation board core1 PLL ratio (cfg_core1_pll)"
    }

    cdl_option CYGHWR_HAL_POWERPC_BUS_SPEED {
        display          "Bus speed (MHz)"
        flavor           data
        default_value    533
        description      "
             MPC8572DS DDRAM bus runs at 533MHz. This is the default setting, with the DDR_CLK
             configured to 66.666MHz and CFG_DDR_PLL set to 8."
    }

    cdl_option CYGHWR_HAL_POWERPC_CPU_CORE_SPEED {
        display          "CPU core (core0) speed (MHz)"
        flavor           data
        calculated       { CYGHWR_HAL_POWERPC_CPU_SPEED * CYGHWR_HAL_POWERPC_MPC8572DS_CORE0_PLL_RATIO }
        description      "
            MPC8572DS core clk runs at 1500MHz. This is the default value, with CCB clock 
            running at 600MHz and CFG_CORE_PLL set to 2.5."
    }

    cdl_option CYGHWR_HAL_POWERPC_CPU_CORE1_SPEED {
        display          "CPU core (core1) speed (MHz)"
        flavor           data
        calculated       { CYGHWR_HAL_POWERPC_CPU_SPEED * CYGHWR_HAL_POWERPC_MPC8572DS_CORE1_PLL_RATIO }
        description      "
            MPC8572DS core1 clk runs at 1500MHz. This is the default value, with CCB clock 
            running at 600MHz and CFG_CORE_PLL set to 2.5."
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        description   "
            Period is bus clock/4/CYGNUM_HAL_RTC_DENOMINATOR."
        flavor        none
        no_define
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
            description   "
              This option selects the number of system clock 'ticks'
              per second.  This rate is sometimes known as the heartbeat rate."
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    { (((CYGHWR_HAL_POWERPC_CPU_SPEED*1000000)/8)/CYGNUM_HAL_RTC_DENOMINATOR) }
        }
    }

    cdl_component CYGPKG_HAL_POWERPC_MPC8572DS_PM {
      display           "Setup performance monitoring on MPC8572DS board"
      default_value     0
      requires          CYGHWR_HAL_POWERPC_ENABLE_PM

      compile plf_pm.c

      description "
                This option allows compilation of performance monitoring example."

      cdl_option CYGSEM_HAL_POWERPC_MPC8572DS_MONITOR_CACHE {
          display       "Monitoring cache operations"
          requires      ! CYGSEM_HAL_POWERPC_MPC8572DS_MONITOR_IO
          default_value 0
          description   "Include/Compile example code for monitoring cache operations."
        }
      cdl_option CYGSEM_HAL_POWERPC_MPC8572DS_MONITOR_IO {
          display       "Monitoring IO operations"
          requires     ! CYGSEM_HAL_POWERPC_MPC8572DS_MONITOR_CACHE
          default_value 0
          description   "Include/Compile example code for monitoring IO operations."
        }
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        description   "
        Global build options including control over
        compiler flags, linker flags and choice of toolchain."

        parent  CYGPKG_NONE

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "powerpc-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { "-msoft-float -mno-hard-dfp -Wa,-me500x2 -Wall -Wpointer-arith -Wstrict-prototypes -Winline -Wundef -Woverloaded-virtual -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc" }
            description   "
                This option controls the global compiler flags which
                are used to compile all packages by
                default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { "-msoft-float -mno-hard-dfp -Wa,-me500x2 -g -nostdlib -Wl,--gc-sections -Wl,-static" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }

        cdl_option CYGBLD_BUILD_GDB_STUBS {
            display "Build GDB stub ROM image"
            default_value 0
            requires { (CYG_HAL_STARTUP == "ROM") || (CYG_HAL_STARTUP == "ROMRAM") }
            requires CYGSEM_HAL_ROM_MONITOR
            requires CYGBLD_BUILD_COMMON_GDB_STUBS
            requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS

            requires CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
            requires CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
            requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
            requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
            no_define
            description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the platform CDL takes care of creating
                an S-Record data file. -- This needs more work"

            make -priority 320 {
                <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
                $(OBJCOPY) -O srec --srec-forceS3 $< $(@:.bin=.s19)
                $(OBJCOPY) -O binary $< $@
            }
        }
    }

    cdl_component CYGPKG_HAL_POWERPC_MPC8572DS_OPTIONS {
        display "MPC8572DS build options"
        flavor  none
        description   "
        Package specific build options including control over
        compiler flags used only in building this package,
        and details of which tests are built."


        cdl_option CYGPKG_HAL_POWERPC_MPC8572DS_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the MPC8572DS HAL. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_HAL_POWERPC_MPC8572DS_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the MPC8572DS HAL. These flags are removed from
                the set of global flags if present."
        }
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM"    ? "powerpc_mpc8572ds_ram" : \
                     CYG_HAL_STARTUP == "ROM"    ? "powerpc_mpc8572ds_rom" : \
                     CYG_HAL_STARTUP == "RAMRAM" ? "powerpc_mpc8572ds_ramram" : \
                                                   "powerpc_mpc8572ds_romram" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM"          ? "<pkgconf/mlt_powerpc_mpc8572ds_ram.ldi>"     : \
                         CYG_HAL_STARTUP == "ROM"          ? "<pkgconf/mlt_powerpc_mpc8572ds_rom.ldi>"     : \
                                                             "<pkgconf/mlt_powerpc_mpc8572ds_romram.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM"          ? "<pkgconf/mlt_powerpc_mpc8572ds_ram.h>"     : \
                         CYG_HAL_STARTUP == "ROM"          ? "<pkgconf/mlt_powerpc_mpc8572ds_rom.h>"     : \
                                                             "<pkgconf/mlt_powerpc_mpc8572ds_romram.h>" }
        }
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { (CYG_HAL_STARTUP == "ROM") || (CYG_HAL_STARTUP == "ROMRAM") }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        bool
        default_value { (CYG_HAL_STARTUP == "RAM" &&
                        !CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS &&
                        !CYGINT_HAL_USE_ROM_MONITOR_UNSUPPORTED &&
                        !CYGSEM_HAL_POWERPC_COPY_VECTORS) ? 1 : 0 }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "RAM" }
        requires      ! CYGSEM_HAL_POWERPC_COPY_VECTORS
        requires      ! CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
        requires      ! CYGINT_HAL_USE_ROM_MONITOR_UNSUPPORTED
        description   "
            Allow coexistence with ROM monitor (CygMon or GDB stubs) by
            only initializing interrupt vectors on startup, thus leaving
            exception handling to the ROM monitor."
    }


    # FIXME: the option above should be adjusted to select between monitor
    #        variants
    cdl_option CYGSEM_HAL_USE_ROM_MONITOR_GDB_stubs {
        parent        CYGPKG_HAL_ROM_MONITOR
        display "Bad CDL workaround"
        calculated 1
        active_if CYGSEM_HAL_USE_ROM_MONITOR
    }


    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGSEM_REDBOOT_PLF_LINUX_BOOT {
            active_if      CYGBLD_BUILD_REDBOOT_WITH_EXEC
            display        "Support booting Linux via RedBoot"
            flavor         bool
            default_value  1
            description    "
               This option enables RedBoot to support booting of a Linux kernel."

            compile plf_redboot_linux_exec.c
        }

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
            image to a binary image suitable for ROM programming.
            This needs more work."

            make -priority 325 {
                <PREFIX>/bin/redboot.bin : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $(@:.bin=.srec)
                $(OBJCOPY) -O binary $< $@
            }
        }
        
        cdl_option CYGHWR_HAL_POWERPC_FORCE_VECTOR_BASE_LOW {
        display          "Force vector base at address 0x0000 0000"
        flavor           bool
        calculated       1
        description      "
             The powerpc architecture allows the vectorbase to live at either
             0x0000 0000 or 0xfff0 0000."
        }
    }
}
