# ==========================================================================
#
#      mini_stm32_fb.cdl
#
#      ILI9325 LCD controller platform specific code
#
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2011 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    ccoutand
# Contributors: 
# Date:         2011-07-01
# Purpose:      
# Description:  ILI9325 LCD controller platform specific code (MINI STM32)
#
#####DESCRIPTIONEND####
#
# ===========================================================================

cdl_package CYGPKG_DEVS_FRAMEBUF_CORTEXM_MINI_STM32 {
    display       "Platform specific device driver for ILI9325 LCD controller (MINI STM32)"
    parent        CYGPKG_DEVS_FRAMEBUF_ILI9325
    active_if     CYGPKG_IO_FRAMEBUF
    active_if     CYGPKG_DEVS_FRAMEBUF_ILI9325
    active_if     CYGPKG_HAL_CORTEXM_STM32

    implements    CYGINT_DEVS_FRAMEBUF_ILI9325_PLF

    include_dir   cyg/io
    compile ili9325_plf.c

    description   "
        This package provides the macros necessary for the ILI9325 
        framebuffer device driver to access the hardware. The ILI9325
        LCD controller initialization sequence is also provided by 
        this package."

    define_proc {
        puts $::cdl_system_header "#define CYGPKG_DEVS_FRAMEBUF_ILI9325_PLF_H <pkgconf/devs_framebuf_cortexm_mini_stm32.h>"
        puts $::cdl_system_header "#define CYGPKG_DEVS_FRAMEBUF_ILI9325_PLF_INL <cyg/io/ili9325_plf.inl>"
    }

    cdl_component CYGPKG_DEVS_FRAMEBUF_CORTEXM_MINI_STM32_OPTIONS {
        display       "Mini STM32 Framebuffer build options"
        flavor        none
        description   "
            Package specific build options including control over
            compiler flags used only in building the generic frame
            buffer package, and details of which tests are built."

        cdl_option CYGPKG_DEVS_FRAMEBUF_CORTEXM_MINI_STM32_TESTS {
            display      "Mini STM32 Framebuffer tests"
            active_if    CYGINT_IO_FRAMEBUF_DEVICES
            flavor       data
            calculated   { "tests/mini_stm32_fb" }
            description "
                This option specifies the set of tests for the Mini STM32 framebuffer package"
        }
    }
}