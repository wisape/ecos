# ==========================================================================
#
#      tsec_eth_drivers.cdl
#
#      Fast ethernet device driver for PowerPC MPC83xx, MPC85xx boards
#
##==========================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 2008 Free Software Foundation, Inc.                        
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
##==========================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):    Edgar Grimberg
# Contributors: ccoutand
# Date:         2009-11-01
# Purpose:      
# Description:  Hardware driver for Freescale eTSEC
#
#####DESCRIPTIONEND####
#
# ===========================================================================

cdl_package CYGPKG_DEVS_ETH_POWERPC_TSEC {
    display       "Freescale PowerQUICC TSEC Ethernet driver"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_POWERPC 
    active_if     CYGPKG_HAL_POWERPC_QUICC2 || CYGPKG_HAL_POWERPC_QUICC3

    include_dir   cyg/io

    description   "Fast ethernet driver for PowerPC MPC83xx/MPC85xx boards."
    compile       -library=libextras.a tsec.c

    # Debug I/O during network stack initialization is not reliable
    # requires { !CYGPKG_NET || CYGPKG_NET_FORCE_SERIAL_CONSOLE == 1 }

    cdl_option CYGNUM_DEVS_ETH_POWERPC_TSEC_BUFSIZE_TX {
        display       "Buffer size"
        flavor        data
        default_value 1536
        description   "
            This option specifies the size of the internal buffers used
            for the PowerPC TSEC/ethernet device."
    }

    cdl_option CYGNUM_DEVS_ETH_POWERPC_TSEC_BUFSIZE_RX {
        display       "Buffer size"
        flavor        data
        default_value 1536
        description   "
            This option specifies the size of the internal buffers used
            for the PowerPC TSEC/ethernet device."
    }

    cdl_option CYGNUM_DEVS_ETH_POWERPC_TSEC_TxNUM {
        display       "Number of output buffers"
        flavor        data
        legal_values  2 to 512
        default_value 64
        description   "
            This option specifies the number of output buffer packets
            to be used for the PowerPC TSEC/ethernet device."
    }

    cdl_option CYGNUM_DEVS_ETH_POWERPC_TSEC_RxNUM {
        display       "Number of input buffers"
        flavor        data
        legal_values  2 to 512
        default_value 64
        description   "
            This option specifies the number of input buffer packets
            to be used for the PowerPC TSEC/ethernet device."
    }

    cdl_option CYGSEM_DEVS_ETH_POWERPC_TSEC_CHATTER {
        display         "Display status messages during Ethernet operations"
        flavor          bool
        default_value   0
        description     "
           Selecting this option will cause the TSEC code to print status
           messages as various Ethernet operations are undertaken."
    }

    cdl_option CYGPKG_DEVS_ETH_POWERPC_TSEC_RMII {
        display         "Reduced-pin mode for 10/100 interfaces"
        flavor          bool
        default_value   0
        description     "
           If this bit is set, a RMII pin interface is expected. Valid only if
           FIFM = 0 and TBIM = 0. RPM and RMM are never set together."
    }

    cdl_component CYGSEM_DEVS_ETH_POWERPC_TSEC_RESET_PHY {
        display       "Reset and reconfigure PHY"
        flavor        bool
        default_value { CYG_HAL_STARTUP != "RAM" }
        active_if     CYGPKG_DEVS_ETH_PHY
        description "
            This option allows control over the physical transceiver"

        cdl_option CYGNUM_DEVS_ETH_POWERPC_TSEC_LINK_MODE {
            display       "Initial link mode"
            flavor        data
            legal_values  { "10Mb" "100Mb" "1000Mb" "Auto" }
            default_value { "Auto" }
            description   "
                This option specifies initial mode for the physical
                link.  The PHY will be reset and then set to this mode."
        }
    }

    cdl_component CYGPKG_DEVS_ETH_POWERPC_TSEC_OPTIONS {
        display "Freescale PowerQUICC TSEC Ethernet driver build options"
        flavor  none
        no_define

        cdl_option CYGPKG_DEVS_ETH_POWERPC_TSEC_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS" }
            description   "
                This option modifies the set of compiler flags for
                building the TSEC ethernet driver package. 
                These flags are used in addition to the set of global 
                flags."
        }
    }

}
